library verilog;
use verilog.vl_types.all;
entity Calculator_tb is
end Calculator_tb;
